`define VEC_SIZE 4
`define VEC_ADDR_WIDTH 3
`define VEC_XPR_LEN (`XPR_LEN * `VEC_SIZE)
