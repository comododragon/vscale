`define XVEC_SIZE 4
`define XVEC_VEC_LEN 29
`define XVEC_NORM_BITS_REM (`XPR_LEN * (`XVEC_VEC_LEN - 1))
`define XVEC_REG_ADDR_WIDTH `REG_ADDR_WIDTH + 1

`define XVEC_OP 7'b0001011
`define XVEC_OP_IMM 7'b0101011
